`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/03/01 16:11:38
// Design Name: 
// Module Name: RGB_Decoder
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module RGB_Decoder(in, out);
    input [2:0] in; // 3��Ʈ�� �Է°��� �޴´�. 
    output reg [5:0] out; // register�� ���� 6��Ʈ�� ��°��� �޴´�. 6��Ʈ�� �޴� ������ LED 2�� �� ���� RGB�� �����Ǿ� �־ ������ ���� ��Ÿ���� �����̴�. 
    
    // Module Body
    always@(*) // always ���� ����Ͽ� ��°��� �Է°��� �����ǰ� �ڵ带 �ۼ��Ѵ�. 
    begin
        case(in)
        // ��찡 �����Ƿ� case���� ���� �ڵ带 �ۼ��Ѵ�.
        3'b000 : out <= 6'b100100; // ���Ǿ��� ����ǥ�� ���� red ���� ��Ÿ���� ���� 6��Ʈ 100100�� out�� �Ҵ��Ѵ�.
        3'b001 : out <= 6'b101101; // ���Ǿ��� ����ǥ�� ���� magenta ���� ��Ÿ���� ���� 6��Ʈ 101101�� out�� �Ҵ��Ѵ�
        3'b010 : out <= 6'b110110; // ���Ǿ��� ����ǥ�� ���� yellow ���� ��Ÿ���� ���� 6��Ʈ 100100�� out�� �Ҵ��Ѵ�
        3'b011 : out <= 6'b010010; // ���Ǿ��� ����ǥ�� ���� green ���� ��Ÿ���� ���� 6��Ʈ 010010�� out�� �Ҵ��Ѵ�
        3'b100 : out <= 6'b011011; // ���Ǿ��� ����ǥ�� ���� cyan ���� ��Ÿ���� ���� 6��Ʈ 011011�� out�� �Ҵ��Ѵ�
        3'b101 : out <= 6'b001001; // ���Ǿ��� ����ǥ�� ���� blue ���� ��Ÿ���� ���� 6��Ʈ 001001�� out�� �Ҵ��Ѵ�
        3'b110 : out <= 6'b111111; // ���Ǿ��� ����ǥ�� ���� white ���� ��Ÿ���� ���� 6��Ʈ 111111�� out�� �Ҵ��Ѵ�
        default : out <= 6'b000000;  // ���� case�� �ش��ϴ� ���� ���� ��� �⺻���� LED off ���� ��Ÿ���� ���� 6��Ʈ 000000�� out�� �Ҵ��Ѵ�
        endcase
    end
endmodule 

